library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sinewavegenerator is
	port(
		clk : in std_logic;
		reset : in std_logic;
		tuningword : in std_logic_vector(7 downto 0);
		sin_out : out std_logic_vector(7 downto 0)
	);
end sinewavegenerator;

architecture rtl of sinewavegenerator is 

    signal phase_acc : unsigned(15 downto 0) := (others => '0');  -- 16-bittinen vaiheakkumulaattori
    signal table_index : unsigned(9 downto 0);                    -- 10-bittinen osoite taulukolle
    signal sin_value : unsigned(7 downto 0);                      -- 8-bittinen siniaallon arvo

	 type t_sin_table is array(0 to 1023) of integer range 0 to 255;
	 constant c_sin_table : t_sin_table := (
		 0 => 127,
		 1 => 128,
		 2 => 129,
		 3 => 129,
		 4 => 130,
		 5 => 131,
		 6 => 132,
		 7 => 132,
		 8 => 133,
		 9 => 134,
		 10 => 135,
		 11 => 136,
		 12 => 136,
		 13 => 137,
		 14 => 138,
		 15 => 139,
		 16 => 139,
		 17 => 140,
		 18 => 141,
		 19 => 142,
		 20 => 143,
		 21 => 143,
		 22 => 144,
		 23 => 145,
		 24 => 146,
		 25 => 146,
		 26 => 147,
		 27 => 148,
		 28 => 149,
		 29 => 150,
		 30 => 150,
		 31 => 151,
		 32 => 152,
		 33 => 153,
		 34 => 153,
		 35 => 154,
		 36 => 155,
		 37 => 156,
		 38 => 156,
		 39 => 157,
		 40 => 158,
		 41 => 159,
		 42 => 159,
		 43 => 160,
		 44 => 161,
		 45 => 162,
		 46 => 163,
		 47 => 163,
		 48 => 164,
		 49 => 165,
		 50 => 166,
		 51 => 166,
		 52 => 167,
		 53 => 168,
		 54 => 168,
		 55 => 169,
		 56 => 170,
		 57 => 171,
		 58 => 171,
		 59 => 172,
		 60 => 173,
		 61 => 174,
		 62 => 174,
		 63 => 175,
		 64 => 176,
		 65 => 177,
		 66 => 177,
		 67 => 178,
		 68 => 179,
		 69 => 179,
		 70 => 180,
		 71 => 181,
		 72 => 182,
		 73 => 182,
		 74 => 183,
		 75 => 184,
		 76 => 184,
		 77 => 185,
		 78 => 186,
		 79 => 186,
		 80 => 187,
		 81 => 188,
		 82 => 188,
		 83 => 189,
		 84 => 190,
		 85 => 191,
		 86 => 191,
		 87 => 192,
		 88 => 193,
		 89 => 193,
		 90 => 194,
		 91 => 195,
		 92 => 195,
		 93 => 196,
		 94 => 197,
		 95 => 197,
		 96 => 198,
		 97 => 198,
		 98 => 199,
		 99 => 200,
		 100 => 200,
		 101 => 201,
		 102 => 202,
		 103 => 202,
		 104 => 203,
		 105 => 204,
		 106 => 204,
		 107 => 205,
		 108 => 205,
		 109 => 206,
		 110 => 207,
		 111 => 207,
		 112 => 208,
		 113 => 208,
		 114 => 209,
		 115 => 210,
		 116 => 210,
		 117 => 211,
		 118 => 211,
		 119 => 212,
		 120 => 213,
		 121 => 213,
		 122 => 214,
		 123 => 214,
		 124 => 215,
		 125 => 215,
		 126 => 216,
		 127 => 217,
		 128 => 217,
		 129 => 218,
		 130 => 218,
		 131 => 219,
		 132 => 219,
		 133 => 220,
		 134 => 220,
		 135 => 221,
		 136 => 221,
		 137 => 222,
		 138 => 223,
		 139 => 223,
		 140 => 224,
		 141 => 224,
		 142 => 225,
		 143 => 225,
		 144 => 226,
		 145 => 226,
		 146 => 227,
		 147 => 227,
		 148 => 228,
		 149 => 228,
		 150 => 228,
		 151 => 229,
		 152 => 229,
		 153 => 230,
		 154 => 230,
		 155 => 231,
		 156 => 231,
		 157 => 232,
		 158 => 232,
		 159 => 233,
		 160 => 233,
		 161 => 233,
		 162 => 234,
		 163 => 234,
		 164 => 235,
		 165 => 235,
		 166 => 236,
		 167 => 236,
		 168 => 236,
		 169 => 237,
		 170 => 237,
		 171 => 238,
		 172 => 238,
		 173 => 238,
		 174 => 239,
		 175 => 239,
		 176 => 239,
		 177 => 240,
		 178 => 240,
		 179 => 241,
		 180 => 241,
		 181 => 241,
		 182 => 242,
		 183 => 242,
		 184 => 242,
		 185 => 243,
		 186 => 243,
		 187 => 243,
		 188 => 244,
		 189 => 244,
		 190 => 244,
		 191 => 244,
		 192 => 245,
		 193 => 245,
		 194 => 245,
		 195 => 246,
		 196 => 246,
		 197 => 246,
		 198 => 247,
		 199 => 247,
		 200 => 247,
		 201 => 247,
		 202 => 248,
		 203 => 248,
		 204 => 248,
		 205 => 248,
		 206 => 249,
		 207 => 249,
		 208 => 249,
		 209 => 249,
		 210 => 249,
		 211 => 250,
		 212 => 250,
		 213 => 250,
		 214 => 250,
		 215 => 250,
		 216 => 251,
		 217 => 251,
		 218 => 251,
		 219 => 251,
		 220 => 251,
		 221 => 252,
		 222 => 252,
		 223 => 252,
		 224 => 252,
		 225 => 252,
		 226 => 252,
		 227 => 252,
		 228 => 253,
		 229 => 253,
		 230 => 253,
		 231 => 253,
		 232 => 253,
		 233 => 253,
		 234 => 253,
		 235 => 253,
		 236 => 254,
		 237 => 254,
		 238 => 254,
		 239 => 254,
		 240 => 254,
		 241 => 254,
		 242 => 254,
		 243 => 254,
		 244 => 254,
		 245 => 254,
		 246 => 254,
		 247 => 254,
		 248 => 254,
		 249 => 254,
		 250 => 254,
		 251 => 254,
		 252 => 254,
		 253 => 254,
		 254 => 254,
		 255 => 254,
		 256 => 255,
		 257 => 254,
		 258 => 254,
		 259 => 254,
		 260 => 254,
		 261 => 254,
		 262 => 254,
		 263 => 254,
		 264 => 254,
		 265 => 254,
		 266 => 254,
		 267 => 254,
		 268 => 254,
		 269 => 254,
		 270 => 254,
		 271 => 254,
		 272 => 254,
		 273 => 254,
		 274 => 254,
		 275 => 254,
		 276 => 254,
		 277 => 253,
		 278 => 253,
		 279 => 253,
		 280 => 253,
		 281 => 253,
		 282 => 253,
		 283 => 253,
		 284 => 253,
		 285 => 252,
		 286 => 252,
		 287 => 252,
		 288 => 252,
		 289 => 252,
		 290 => 252,
		 291 => 252,
		 292 => 251,
		 293 => 251,
		 294 => 251,
		 295 => 251,
		 296 => 251,
		 297 => 250,
		 298 => 250,
		 299 => 250,
		 300 => 250,
		 301 => 250,
		 302 => 249,
		 303 => 249,
		 304 => 249,
		 305 => 249,
		 306 => 249,
		 307 => 248,
		 308 => 248,
		 309 => 248,
		 310 => 248,
		 311 => 247,
		 312 => 247,
		 313 => 247,
		 314 => 247,
		 315 => 246,
		 316 => 246,
		 317 => 246,
		 318 => 245,
		 319 => 245,
		 320 => 245,
		 321 => 244,
		 322 => 244,
		 323 => 244,
		 324 => 244,
		 325 => 243,
		 326 => 243,
		 327 => 243,
		 328 => 242,
		 329 => 242,
		 330 => 242,
		 331 => 241,
		 332 => 241,
		 333 => 241,
		 334 => 240,
		 335 => 240,
		 336 => 239,
		 337 => 239,
		 338 => 239,
		 339 => 238,
		 340 => 238,
		 341 => 238,
		 342 => 237,
		 343 => 237,
		 344 => 236,
		 345 => 236,
		 346 => 236,
		 347 => 235,
		 348 => 235,
		 349 => 234,
		 350 => 234,
		 351 => 233,
		 352 => 233,
		 353 => 233,
		 354 => 232,
		 355 => 232,
		 356 => 231,
		 357 => 231,
		 358 => 230,
		 359 => 230,
		 360 => 229,
		 361 => 229,
		 362 => 228,
		 363 => 228,
		 364 => 228,
		 365 => 227,
		 366 => 227,
		 367 => 226,
		 368 => 226,
		 369 => 225,
		 370 => 225,
		 371 => 224,
		 372 => 224,
		 373 => 223,
		 374 => 223,
		 375 => 222,
		 376 => 221,
		 377 => 221,
		 378 => 220,
		 379 => 220,
		 380 => 219,
		 381 => 219,
		 382 => 218,
		 383 => 218,
		 384 => 217,
		 385 => 217,
		 386 => 216,
		 387 => 215,
		 388 => 215,
		 389 => 214,
		 390 => 214,
		 391 => 213,
		 392 => 213,
		 393 => 212,
		 394 => 211,
		 395 => 211,
		 396 => 210,
		 397 => 210,
		 398 => 209,
		 399 => 208,
		 400 => 208,
		 401 => 207,
		 402 => 207,
		 403 => 206,
		 404 => 205,
		 405 => 205,
		 406 => 204,
		 407 => 204,
		 408 => 203,
		 409 => 202,
		 410 => 202,
		 411 => 201,
		 412 => 200,
		 413 => 200,
		 414 => 199,
		 415 => 198,
		 416 => 198,
		 417 => 197,
		 418 => 197,
		 419 => 196,
		 420 => 195,
		 421 => 195,
		 422 => 194,
		 423 => 193,
		 424 => 193,
		 425 => 192,
		 426 => 191,
		 427 => 191,
		 428 => 190,
		 429 => 189,
		 430 => 188,
		 431 => 188,
		 432 => 187,
		 433 => 186,
		 434 => 186,
		 435 => 185,
		 436 => 184,
		 437 => 184,
		 438 => 183,
		 439 => 182,
		 440 => 182,
		 441 => 181,
		 442 => 180,
		 443 => 179,
		 444 => 179,
		 445 => 178,
		 446 => 177,
		 447 => 177,
		 448 => 176,
		 449 => 175,
		 450 => 174,
		 451 => 174,
		 452 => 173,
		 453 => 172,
		 454 => 171,
		 455 => 171,
		 456 => 170,
		 457 => 169,
		 458 => 168,
		 459 => 168,
		 460 => 167,
		 461 => 166,
		 462 => 166,
		 463 => 165,
		 464 => 164,
		 465 => 163,
		 466 => 163,
		 467 => 162,
		 468 => 161,
		 469 => 160,
		 470 => 159,
		 471 => 159,
		 472 => 158,
		 473 => 157,
		 474 => 156,
		 475 => 156,
		 476 => 155,
		 477 => 154,
		 478 => 153,
		 479 => 153,
		 480 => 152,
		 481 => 151,
		 482 => 150,
		 483 => 150,
		 484 => 149,
		 485 => 148,
		 486 => 147,
		 487 => 146,
		 488 => 146,
		 489 => 145,
		 490 => 144,
		 491 => 143,
		 492 => 143,
		 493 => 142,
		 494 => 141,
		 495 => 140,
		 496 => 139,
		 497 => 139,
		 498 => 138,
		 499 => 137,
		 500 => 136,
		 501 => 136,
		 502 => 135,
		 503 => 134,
		 504 => 133,
		 505 => 132,
		 506 => 132,
		 507 => 131,
		 508 => 130,
		 509 => 129,
		 510 => 129,
		 511 => 128,
		 512 => 127,
		 513 => 126,
		 514 => 125,
		 515 => 125,
		 516 => 124,
		 517 => 123,
		 518 => 122,
		 519 => 122,
		 520 => 121,
		 521 => 120,
		 522 => 119,
		 523 => 118,
		 524 => 118,
		 525 => 117,
		 526 => 116,
		 527 => 115,
		 528 => 115,
		 529 => 114,
		 530 => 113,
		 531 => 112,
		 532 => 111,
		 533 => 111,
		 534 => 110,
		 535 => 109,
		 536 => 108,
		 537 => 108,
		 538 => 107,
		 539 => 106,
		 540 => 105,
		 541 => 104,
		 542 => 104,
		 543 => 103,
		 544 => 102,
		 545 => 101,
		 546 => 101,
		 547 => 100,
		 548 => 99,
		 549 => 98,
		 550 => 98,
		 551 => 97,
		 552 => 96,
		 553 => 95,
		 554 => 95,
		 555 => 94,
		 556 => 93,
		 557 => 92,
		 558 => 91,
		 559 => 91,
		 560 => 90,
		 561 => 89,
		 562 => 88,
		 563 => 88,
		 564 => 87,
		 565 => 86,
		 566 => 86,
		 567 => 85,
		 568 => 84,
		 569 => 83,
		 570 => 83,
		 571 => 82,
		 572 => 81,
		 573 => 80,
		 574 => 80,
		 575 => 79,
		 576 => 78,
		 577 => 77,
		 578 => 77,
		 579 => 76,
		 580 => 75,
		 581 => 75,
		 582 => 74,
		 583 => 73,
		 584 => 72,
		 585 => 72,
		 586 => 71,
		 587 => 70,
		 588 => 70,
		 589 => 69,
		 590 => 68,
		 591 => 68,
		 592 => 67,
		 593 => 66,
		 594 => 66,
		 595 => 65,
		 596 => 64,
		 597 => 63,
		 598 => 63,
		 599 => 62,
		 600 => 61,
		 601 => 61,
		 602 => 60,
		 603 => 59,
		 604 => 59,
		 605 => 58,
		 606 => 57,
		 607 => 57,
		 608 => 56,
		 609 => 56,
		 610 => 55,
		 611 => 54,
		 612 => 54,
		 613 => 53,
		 614 => 52,
		 615 => 52,
		 616 => 51,
		 617 => 50,
		 618 => 50,
		 619 => 49,
		 620 => 49,
		 621 => 48,
		 622 => 47,
		 623 => 47,
		 624 => 46,
		 625 => 46,
		 626 => 45,
		 627 => 44,
		 628 => 44,
		 629 => 43,
		 630 => 43,
		 631 => 42,
		 632 => 41,
		 633 => 41,
		 634 => 40,
		 635 => 40,
		 636 => 39,
		 637 => 39,
		 638 => 38,
		 639 => 37,
		 640 => 37,
		 641 => 36,
		 642 => 36,
		 643 => 35,
		 644 => 35,
		 645 => 34,
		 646 => 34,
		 647 => 33,
		 648 => 33,
		 649 => 32,
		 650 => 31,
		 651 => 31,
		 652 => 30,
		 653 => 30,
		 654 => 29,
		 655 => 29,
		 656 => 28,
		 657 => 28,
		 658 => 27,
		 659 => 27,
		 660 => 26,
		 661 => 26,
		 662 => 26,
		 663 => 25,
		 664 => 25,
		 665 => 24,
		 666 => 24,
		 667 => 23,
		 668 => 23,
		 669 => 22,
		 670 => 22,
		 671 => 21,
		 672 => 21,
		 673 => 21,
		 674 => 20,
		 675 => 20,
		 676 => 19,
		 677 => 19,
		 678 => 18,
		 679 => 18,
		 680 => 18,
		 681 => 17,
		 682 => 17,
		 683 => 16,
		 684 => 16,
		 685 => 16,
		 686 => 15,
		 687 => 15,
		 688 => 15,
		 689 => 14,
		 690 => 14,
		 691 => 13,
		 692 => 13,
		 693 => 13,
		 694 => 12,
		 695 => 12,
		 696 => 12,
		 697 => 11,
		 698 => 11,
		 699 => 11,
		 700 => 10,
		 701 => 10,
		 702 => 10,
		 703 => 10,
		 704 => 9,
		 705 => 9,
		 706 => 9,
		 707 => 8,
		 708 => 8,
		 709 => 8,
		 710 => 7,
		 711 => 7,
		 712 => 7,
		 713 => 7,
		 714 => 6,
		 715 => 6,
		 716 => 6,
		 717 => 6,
		 718 => 5,
		 719 => 5,
		 720 => 5,
		 721 => 5,
		 722 => 5,
		 723 => 4,
		 724 => 4,
		 725 => 4,
		 726 => 4,
		 727 => 4,
		 728 => 3,
		 729 => 3,
		 730 => 3,
		 731 => 3,
		 732 => 3,
		 733 => 2,
		 734 => 2,
		 735 => 2,
		 736 => 2,
		 737 => 2,
		 738 => 2,
		 739 => 2,
		 740 => 1,
		 741 => 1,
		 742 => 1,
		 743 => 1,
		 744 => 1,
		 745 => 1,
		 746 => 1,
		 747 => 1,
		 748 => 0,
		 749 => 0,
		 750 => 0,
		 751 => 0,
		 752 => 0,
		 753 => 0,
		 754 => 0,
		 755 => 0,
		 756 => 0,
		 757 => 0,
		 758 => 0,
		 759 => 0,
		 760 => 0,
		 761 => 0,
		 762 => 0,
		 763 => 0,
		 764 => 0,
		 765 => 0,
		 766 => 0,
		 767 => 0,
		 768 => 0,
		 769 => 0,
		 770 => 0,
		 771 => 0,
		 772 => 0,
		 773 => 0,
		 774 => 0,
		 775 => 0,
		 776 => 0,
		 777 => 0,
		 778 => 0,
		 779 => 0,
		 780 => 0,
		 781 => 0,
		 782 => 0,
		 783 => 0,
		 784 => 0,
		 785 => 0,
		 786 => 0,
		 787 => 0,
		 788 => 0,
		 789 => 1,
		 790 => 1,
		 791 => 1,
		 792 => 1,
		 793 => 1,
		 794 => 1,
		 795 => 1,
		 796 => 1,
		 797 => 2,
		 798 => 2,
		 799 => 2,
		 800 => 2,
		 801 => 2,
		 802 => 2,
		 803 => 2,
		 804 => 3,
		 805 => 3,
		 806 => 3,
		 807 => 3,
		 808 => 3,
		 809 => 4,
		 810 => 4,
		 811 => 4,
		 812 => 4,
		 813 => 4,
		 814 => 5,
		 815 => 5,
		 816 => 5,
		 817 => 5,
		 818 => 5,
		 819 => 6,
		 820 => 6,
		 821 => 6,
		 822 => 6,
		 823 => 7,
		 824 => 7,
		 825 => 7,
		 826 => 7,
		 827 => 8,
		 828 => 8,
		 829 => 8,
		 830 => 9,
		 831 => 9,
		 832 => 9,
		 833 => 10,
		 834 => 10,
		 835 => 10,
		 836 => 10,
		 837 => 11,
		 838 => 11,
		 839 => 11,
		 840 => 12,
		 841 => 12,
		 842 => 12,
		 843 => 13,
		 844 => 13,
		 845 => 13,
		 846 => 14,
		 847 => 14,
		 848 => 15,
		 849 => 15,
		 850 => 15,
		 851 => 16,
		 852 => 16,
		 853 => 16,
		 854 => 17,
		 855 => 17,
		 856 => 18,
		 857 => 18,
		 858 => 18,
		 859 => 19,
		 860 => 19,
		 861 => 20,
		 862 => 20,
		 863 => 21,
		 864 => 21,
		 865 => 21,
		 866 => 22,
		 867 => 22,
		 868 => 23,
		 869 => 23,
		 870 => 24,
		 871 => 24,
		 872 => 25,
		 873 => 25,
		 874 => 26,
		 875 => 26,
		 876 => 26,
		 877 => 27,
		 878 => 27,
		 879 => 28,
		 880 => 28,
		 881 => 29,
		 882 => 29,
		 883 => 30,
		 884 => 30,
		 885 => 31,
		 886 => 31,
		 887 => 32,
		 888 => 33,
		 889 => 33,
		 890 => 34,
		 891 => 34,
		 892 => 35,
		 893 => 35,
		 894 => 36,
		 895 => 36,
		 896 => 37,
		 897 => 37,
		 898 => 38,
		 899 => 39,
		 900 => 39,
		 901 => 40,
		 902 => 40,
		 903 => 41,
		 904 => 41,
		 905 => 42,
		 906 => 43,
		 907 => 43,
		 908 => 44,
		 909 => 44,
		 910 => 45,
		 911 => 46,
		 912 => 46,
		 913 => 47,
		 914 => 47,
		 915 => 48,
		 916 => 49,
		 917 => 49,
		 918 => 50,
		 919 => 50,
		 920 => 51,
		 921 => 52,
		 922 => 52,
		 923 => 53,
		 924 => 54,
		 925 => 54,
		 926 => 55,
		 927 => 56,
		 928 => 56,
		 929 => 57,
		 930 => 57,
		 931 => 58,
		 932 => 59,
		 933 => 59,
		 934 => 60,
		 935 => 61,
		 936 => 61,
		 937 => 62,
		 938 => 63,
		 939 => 63,
		 940 => 64,
		 941 => 65,
		 942 => 66,
		 943 => 66,
		 944 => 67,
		 945 => 68,
		 946 => 68,
		 947 => 69,
		 948 => 70,
		 949 => 70,
		 950 => 71,
		 951 => 72,
		 952 => 72,
		 953 => 73,
		 954 => 74,
		 955 => 75,
		 956 => 75,
		 957 => 76,
		 958 => 77,
		 959 => 77,
		 960 => 78,
		 961 => 79,
		 962 => 80,
		 963 => 80,
		 964 => 81,
		 965 => 82,
		 966 => 83,
		 967 => 83,
		 968 => 84,
		 969 => 85,
		 970 => 86,
		 971 => 86,
		 972 => 87,
		 973 => 88,
		 974 => 88,
		 975 => 89,
		 976 => 90,
		 977 => 91,
		 978 => 91,
		 979 => 92,
		 980 => 93,
		 981 => 94,
		 982 => 95,
		 983 => 95,
		 984 => 96,
		 985 => 97,
		 986 => 98,
		 987 => 98,
		 988 => 99,
		 989 => 100,
		 990 => 101,
		 991 => 101,
		 992 => 102,
		 993 => 103,
		 994 => 104,
		 995 => 104,
		 996 => 105,
		 997 => 106,
		 998 => 107,
		 999 => 108,
		 1000 => 108,
		 1001 => 109,
		 1002 => 110,
		 1003 => 111,
		 1004 => 111,
		 1005 => 112,
		 1006 => 113,
		 1007 => 114,
		 1008 => 115,
		 1009 => 115,
		 1010 => 116,
		 1011 => 117,
		 1012 => 118,
		 1013 => 118,
		 1014 => 119,
		 1015 => 120,
		 1016 => 121,
		 1017 => 122,
		 1018 => 122,
		 1019 => 123,
		 1020 => 124,
		 1021 => 125,
		 1022 => 125,
		 1023 => 126
	);
	 
begin

    -- Prosessi, joka päivittää vaiheakkumulaattorin ja laskee siniaallon
    process(clk)
    begin
        if rising_edge(clk) then
            if reset = '1' then
                phase_acc <= (others => '0');  -- Nollaa vaiheakkumulaattori resetissä
            else
                -- Lisää taajuusohjausluku vaiheakkumulaattoriin (DDS-periaate)
                phase_acc <= phase_acc + unsigned(tuningword & "00000000"); 
            end if;
        end if;
    end process;

    -- Käytä vaiheakkumulaattorin 10 ylimmäistä bittiä taulukon osoitteena
    table_index <= phase_acc(15 downto 6);  -- Osoita siniaaltotaulukkoa

    -- Lue taulukosta siniaallon arvo
    sin_value <= to_unsigned(c_sin_table(to_integer(table_index)), 8);

    -- Lähetä siniaallon arvo ulos 8-bittisenä signaalina
    sin_out <= std_logic_vector(sin_value);


end rtl;